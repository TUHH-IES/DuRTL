module ift_tag_test(a, b, c, d, e);
 input a,b,c,d;
 output e;

 assign e = a & b & c & e;
endmodule

