module split( a, b, out);

	input [5:0] a;
	input [5:0] b;
	output [5:0] out;
	wire [5:0] out;
	integer i;

	assign out = a & i;



endmodule
