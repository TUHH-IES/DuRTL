module d1(a,b);

input a;
output wire b;

assign b = a;

endmodule
