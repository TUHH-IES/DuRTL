module openMSP430( cpu_en, dbg_en, dbg_i2c_addr, dbg_i2c_broadcast, dbg_i2c_scl, dbg_i2c_sda_in, dbg_uart_rxd, dco_clk, dma_addr, dma_din, dma_en, dma_priority, dma_we, dma_wkup, dmem_dout, irq, lfxt_clk, nmi, per_dout, pmem_dout, reset_n, scan_enable, scan_mode, wkup, aclk, aclk_en, dbg_freeze, dbg_i2c_sda_out, dbg_uart_txd, dco_enable, dco_wkup, dma_dout, dma_ready, dma_resp, dmem_addr, dmem_cen, dmem_din, dmem_wen, irq_acc, lfxt_enable, lfxt_wkup, mclk, per_addr, per_din, per_en, per_we, pmem_addr, pmem_cen, pmem_din, pmem_wen, puc_rst, smclk, smclk_en);
input cpu_en;
input dbg_en;
input [6:0] dbg_i2c_addr;
input [6:0] dbg_i2c_broadcast;
input dbg_i2c_scl;
input dbg_i2c_sda_in;
input dbg_uart_rxd;
input dco_clk;
input [14:0] dma_addr;
input [15:0] dma_din;
input dma_en;
input dma_priority;
input [1:0] dma_we;
input dma_wkup;
input [15:0] dmem_dout;
input [13:0] irq;
input lfxt_clk;
input nmi;
input [15:0] per_dout;
input [15:0] pmem_dout;
input reset_n;
input scan_enable;
input scan_mode;
input wkup;
output aclk;
output aclk_en;
output dbg_freeze;
output dbg_i2c_sda_out;
output dbg_uart_txd;
output dco_enable;
output dco_wkup;
output [15:0] dma_dout;
output dma_ready;
output dma_resp;
output [8:0] dmem_addr;
output dmem_cen;
output [15:0] dmem_din;
output [1:0] dmem_wen;
output [13:0] irq_acc;
output lfxt_enable;
output lfxt_wkup;
output mclk;
output [13:0] per_addr;
output [15:0] per_din;
output per_en;
output [1:0] per_we;
output [10:0] pmem_addr;
output pmem_cen;
output [15:0] pmem_din;
output [1:0] pmem_wen;
output puc_rst;
output smclk;
output smclk_en;
m_19 ins( cpu_en, dbg_en, dbg_i2c_addr, dbg_i2c_broadcast, dbg_i2c_scl, dbg_i2c_sda_in, dbg_uart_rxd, dco_clk, dma_addr, dma_din, dma_en, dma_priority, dma_we, dma_wkup, dmem_dout, irq, lfxt_clk, nmi, per_dout, pmem_dout, reset_n, scan_enable, scan_mode, wkup, aclk, aclk_en, dbg_freeze, dbg_i2c_sda_out, dbg_uart_txd, dco_enable, dco_wkup, dma_dout, dma_ready, dma_resp, dmem_addr, dmem_cen, dmem_din, dmem_wen, irq_acc, lfxt_enable, lfxt_wkup, dma_mclk, per_addr, per_din, per_en, per_we, pmem_addr, pmem_cen, pmem_din, pmem_wen, puc_rst, smclk, smclk_en);
endmodule