`timescale 1us/100ns
module tb_pmux_ue();
	reg [1:0] A;
	reg [5:0] B;
	reg [2:0] S;
	wire[1:0] Y;
	

	m_0 d1(.A(A),.B(B),.S(S),.Y(Y));

	initial begin 
		#5;
		 A <= 0;
		 B <= 0;
		 S <= 0;
		 #5;
		 A <= 0;
		 B <= 0;
		 S <= 1;
		 #5;
		 A <= 0;
		 B <= 0;
		 S <= 2;
		 #5;
		 A <= 0;
		 B <= 0;
		 S <= 3;
		 #5;
		 A <= 0;
		 B <= 0;
		 S <= 4;
		 #5;
		 A <= 0;
		 B <= 0;
		 S <= 5;
		 #5;
		 A <= 0;
		 B <= 0;
		 S <= 6;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 0;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 1;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 2;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 3;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 4;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 5;
		 #5;
		 A <= 0;
		 B <= 19;
		 S <= 6;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 0;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 1;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 2;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 3;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 4;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 5;
		 #5;
		 A <= 0;
		 B <= 38;
		 S <= 6;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 0;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 1;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 2;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 3;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 4;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 5;
		 #5;
		 A <= 0;
		 B <= 57;
		 S <= 6;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 0;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 1;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 2;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 3;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 4;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 5;
		 #5;
		 A <= 1;
		 B <= 0;
		 S <= 6;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 0;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 1;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 2;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 3;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 4;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 5;
		 #5;
		 A <= 1;
		 B <= 19;
		 S <= 6;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 0;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 1;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 2;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 3;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 4;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 5;
		 #5;
		 A <= 1;
		 B <= 38;
		 S <= 6;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 0;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 1;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 2;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 3;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 4;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 5;
		 #5;
		 A <= 1;
		 B <= 57;
		 S <= 6;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 0;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 1;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 2;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 3;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 4;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 5;
		 #5;
		 A <= 2;
		 B <= 0;
		 S <= 6;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 0;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 1;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 2;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 3;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 4;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 5;
		 #5;
		 A <= 2;
		 B <= 19;
		 S <= 6;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 0;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 1;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 2;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 3;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 4;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 5;
		 #5;
		 A <= 2;
		 B <= 38;
		 S <= 6;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 0;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 1;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 2;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 3;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 4;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 5;
		 #5;
		 A <= 2;
		 B <= 57;
		 S <= 6;

		 $finish;
	end
	initial
	begin
		$dumpfile(`DUMP_FILE_NAME);
		//$dumpfile("pmux_ue.vcd");
		$dumpvars(1);		//writing the vcd file
	end
 	
endmodule 

