module xorGate( a, b, out);

	input a, b;
	output out;
	wire out;

	assign out = a ^ b;

endmodule
