module M50 (in_0,in_1,out_0,out_1);
   input [16:0] in_0;
   input [16:0] in_1;
   output [16:0] out_0;
   output [16:0] out_1;

   assign out_0 = in_0&in_1;
   assign out_1 = in_0|in_1;
endmodule



module M49 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M50 m0(in_0,in_1,in_2,in_3,in_4,in_5,in_6,in_7,in_8,in_9,in_10,in_11,in_12,in_13,in_14,in_15,in_16,in_17,in_18,in_19,in_20,in_21,in_22,in_23,in_24,in_25,in_26,in_27,in_28,in_29,in_30,in_31,in_32,in_33,in_34,in_35,in_36,in_37,in_38,in_39,in_40,in_41,in_42,in_43,in_44,in_45,in_46,in_47,in_48,w_0,w_1);
   M50 m1(in_49,in_50,in_51,in_52,in_53,in_54,in_55,in_56,in_57,in_58,in_59,in_60,in_61,in_62,in_63,in_64,in_65,in_66,in_67,in_68,in_69,in_70,in_71,in_72,in_73,in_74,in_75,in_76,in_77,in_78,in_79,in_80,in_81,in_82,in_83,in_84,in_85,in_86,in_87,in_88,in_89,in_90,in_91,in_92,in_93,in_94,in_95,in_96,in_97,w_2,w_3);
   M50 m2(in_98,in_99,in_100,in_101,in_102,in_103,in_104,in_105,in_106,in_107,in_108,in_109,in_110,in_111,in_112,in_113,in_114,in_115,in_116,in_117,in_118,in_119,in_120,in_121,in_122,in_123,in_124,in_125,in_126,in_127,in_128,in_129,in_130,in_131,in_132,in_133,in_134,in_135,in_136,in_137,in_138,in_139,in_140,in_141,in_142,in_143,in_144,in_145,in_146,w_4,w_5);
   M50 m3(in_147,in_148,in_149,in_150,in_151,in_152,in_153,in_154,in_155,in_156,in_157,in_158,in_159,in_160,in_161,in_162,in_163,in_164,in_165,in_166,in_167,in_168,in_169,in_170,in_171,in_172,in_173,in_174,in_175,in_176,in_177,in_178,in_179,in_180,in_181,in_182,in_183,in_184,in_185,in_186,in_187,in_188,in_189,in_190,in_191,in_192,in_193,in_194,in_195,w_6,w_7);
   M50 m4(in_196,in_197,in_198,in_199,in_200,in_201,in_202,in_203,in_204,in_205,in_206,in_207,in_208,in_209,in_210,in_211,in_212,in_213,in_214,in_215,in_216,in_217,in_218,in_219,in_220,in_221,in_222,in_223,in_224,in_225,in_226,in_227,in_228,in_229,in_230,in_231,in_232,in_233,in_234,in_235,in_236,in_237,in_238,in_239,in_240,in_241,in_242,in_243,in_244,w_8,w_9);
   M50 m5(in_245,in_246,in_247,in_248,in_249,in_250,in_251,in_252,in_253,in_254,in_255,in_256,in_257,in_258,in_259,in_260,in_261,in_262,in_263,in_264,in_265,in_266,in_267,in_268,in_269,in_270,in_271,in_272,in_273,in_274,in_275,in_276,in_277,in_278,in_279,in_280,in_281,in_282,in_283,in_284,in_285,in_286,in_287,in_288,in_289,in_290,in_291,in_292,in_293,w_10,w_11);
   M50 m6(in_294,in_295,in_296,in_297,in_298,in_299,in_300,in_301,in_302,in_303,in_304,in_305,in_306,in_307,in_308,in_309,in_310,in_311,in_312,in_313,in_314,in_315,in_316,in_317,in_318,in_319,in_320,in_321,in_322,in_323,in_324,in_325,in_326,in_327,in_328,in_329,in_330,in_331,in_332,in_333,in_334,in_335,in_336,in_337,in_338,in_339,in_340,in_341,in_342,w_12,w_13);
   M50 m7(in_343,in_344,in_345,in_346,in_347,in_348,in_349,in_350,in_351,in_352,in_353,in_354,in_355,in_356,in_357,in_358,in_359,in_360,in_361,in_362,in_363,in_364,in_365,in_366,in_367,in_368,in_369,in_370,in_371,in_372,in_373,in_374,in_375,in_376,in_377,in_378,in_379,in_380,in_381,in_382,in_383,in_384,in_385,in_386,in_387,in_388,in_389,in_390,in_391,w_14,w_15);
   M50 m8(in_392,in_393,in_394,in_395,in_396,in_397,in_398,in_399,in_400,in_401,in_402,in_403,in_404,in_405,in_406,in_407,in_408,in_409,in_410,in_411,in_412,in_413,in_414,in_415,in_416,in_417,in_418,in_419,in_420,in_421,in_422,in_423,in_424,in_425,in_426,in_427,in_428,in_429,in_430,in_431,in_432,in_433,in_434,in_435,in_436,in_437,in_438,in_439,in_440,w_16,w_17);
   M50 m9(in_441,in_442,in_443,in_444,in_445,in_446,in_447,in_448,in_449,in_450,in_451,in_452,in_453,in_454,in_455,in_456,in_457,in_458,in_459,in_460,in_461,in_462,in_463,in_464,in_465,in_466,in_467,in_468,in_469,in_470,in_471,in_472,in_473,in_474,in_475,in_476,in_477,in_478,in_479,in_480,in_481,in_482,in_483,in_484,in_485,in_486,in_487,in_488,in_489,w_18,w_19);
   M50 m10(in_490,in_491,in_492,in_493,in_494,in_495,in_496,in_497,in_498,in_499,in_500,in_501,in_502,in_503,in_504,in_505,in_506,in_507,in_508,in_509,in_510,in_511,in_512,in_513,in_514,in_515,in_516,in_517,in_518,in_519,in_520,in_521,in_522,in_523,in_524,in_525,in_526,in_527,in_528,in_529,in_530,in_531,in_532,in_533,in_534,in_535,in_536,in_537,in_538,w_20,w_21);
   M50 m11(in_539,in_540,in_541,in_542,in_543,in_544,in_545,in_546,in_547,in_548,in_549,in_550,in_551,in_552,in_553,in_554,in_555,in_556,in_557,in_558,in_559,in_560,in_561,in_562,in_563,in_564,in_565,in_566,in_567,in_568,in_569,in_570,in_571,in_572,in_573,in_574,in_575,in_576,in_577,in_578,in_579,in_580,in_581,in_582,in_583,in_584,in_585,in_586,in_587,w_22,w_23);
   M50 m12(in_588,in_589,in_590,in_591,in_592,in_593,in_594,in_595,in_596,in_597,in_598,in_599,in_600,in_601,in_602,in_603,in_604,in_605,in_606,in_607,in_608,in_609,in_610,in_611,in_612,in_613,in_614,in_615,in_616,in_617,in_618,in_619,in_620,in_621,in_622,in_623,in_624,in_625,in_626,in_627,in_628,in_629,in_630,in_631,in_632,in_633,in_634,in_635,in_636,w_24,w_25);
   M50 m13(in_637,in_638,in_639,in_640,in_641,in_642,in_643,in_644,in_645,in_646,in_647,in_648,in_649,in_650,in_651,in_652,in_653,in_654,in_655,in_656,in_657,in_658,in_659,in_660,in_661,in_662,in_663,in_664,in_665,in_666,in_667,in_668,in_669,in_670,in_671,in_672,in_673,in_674,in_675,in_676,in_677,in_678,in_679,in_680,in_681,in_682,in_683,in_684,in_685,w_26,w_27);
   M50 m14(in_686,in_687,in_688,in_689,in_690,in_691,in_692,in_693,in_694,in_695,in_696,in_697,in_698,in_699,in_700,in_701,in_702,in_703,in_704,in_705,in_706,in_707,in_708,in_709,in_710,in_711,in_712,in_713,in_714,in_715,in_716,in_717,in_718,in_719,in_720,in_721,in_722,in_723,in_724,in_725,in_726,in_727,in_728,in_729,in_730,in_731,in_732,in_733,in_734,w_28,w_29);
   M50 m15(in_735,in_736,in_737,in_738,in_739,in_740,in_741,in_742,in_743,in_744,in_745,in_746,in_747,in_748,in_749,in_750,in_751,in_752,in_753,in_754,in_755,in_756,in_757,in_758,in_759,in_760,in_761,in_762,in_763,in_764,in_765,in_766,in_767,in_768,in_769,in_770,in_771,in_772,in_773,in_774,in_775,in_776,in_777,in_778,in_779,in_780,in_781,in_782,in_783,w_30,w_31);
   M50 m16(in_784,in_785,in_786,in_787,in_788,in_789,in_790,in_791,in_792,in_793,in_794,in_795,in_796,in_797,in_798,in_799,in_800,in_801,in_802,in_803,in_804,in_805,in_806,in_807,in_808,in_809,in_810,in_811,in_812,in_813,in_814,in_815,in_816,in_817,in_818,in_819,in_820,in_821,in_822,in_823,in_824,in_825,in_826,in_827,in_828,in_829,in_830,in_831,in_832,w_32,w_33);
   M50 m17(in_833,in_834,in_835,in_836,in_837,in_838,in_839,in_840,in_841,in_842,in_843,in_844,in_845,in_846,in_847,in_848,in_849,in_850,in_851,in_852,in_853,in_854,in_855,in_856,in_857,in_858,in_859,in_860,in_861,in_862,in_863,in_864,in_865,in_866,in_867,in_868,in_869,in_870,in_871,in_872,in_873,in_874,in_875,in_876,in_877,in_878,in_879,in_880,in_881,w_34,w_35);
   M50 m18(in_882,in_883,in_884,in_885,in_886,in_887,in_888,in_889,in_890,in_891,in_892,in_893,in_894,in_895,in_896,in_897,in_898,in_899,in_900,in_901,in_902,in_903,in_904,in_905,in_906,in_907,in_908,in_909,in_910,in_911,in_912,in_913,in_914,in_915,in_916,in_917,in_918,in_919,in_920,in_921,in_922,in_923,in_924,in_925,in_926,in_927,in_928,in_929,in_930,w_36,w_37);
   M50 m19(in_931,in_932,in_933,in_934,in_935,in_936,in_937,in_938,in_939,in_940,in_941,in_942,in_943,in_944,in_945,in_946,in_947,in_948,in_949,in_950,in_951,in_952,in_953,in_954,in_955,in_956,in_957,in_958,in_959,in_960,in_961,in_962,in_963,in_964,in_965,in_966,in_967,in_968,in_969,in_970,in_971,in_972,in_973,in_974,in_975,in_976,in_977,in_978,in_979,w_38,w_39);
   M50 m20(in_980,in_981,in_982,in_983,in_984,in_985,in_986,in_987,in_988,in_989,in_990,in_991,in_992,in_993,in_994,in_995,in_996,in_997,in_998,in_999,in_1000,in_1001,in_1002,in_1003,in_1004,in_1005,in_1006,in_1007,in_1008,in_1009,in_1010,in_1011,in_1012,in_1013,in_1014,in_1015,in_1016,in_1017,in_1018,in_1019,in_1020,in_1021,in_1022,in_1023,in_1024,in_1025,in_1026,in_1027,in_1028,w_40,w_41);
   M50 m21(in_1029,in_1030,in_1031,in_1032,in_1033,in_1034,in_1035,in_1036,in_1037,in_1038,in_1039,in_1040,in_1041,in_1042,in_1043,in_1044,in_1045,in_1046,in_1047,in_1048,in_1049,in_1050,in_1051,in_1052,in_1053,in_1054,in_1055,in_1056,in_1057,in_1058,in_1059,in_1060,in_1061,in_1062,in_1063,in_1064,in_1065,in_1066,in_1067,in_1068,in_1069,in_1070,in_1071,in_1072,in_1073,in_1074,in_1075,in_1076,in_1077,w_42,w_43);
   M50 m22(in_1078,in_1079,in_1080,in_1081,in_1082,in_1083,in_1084,in_1085,in_1086,in_1087,in_1088,in_1089,in_1090,in_1091,in_1092,in_1093,in_1094,in_1095,in_1096,in_1097,in_1098,in_1099,in_1100,in_1101,in_1102,in_1103,in_1104,in_1105,in_1106,in_1107,in_1108,in_1109,in_1110,in_1111,in_1112,in_1113,in_1114,in_1115,in_1116,in_1117,in_1118,in_1119,in_1120,in_1121,in_1122,in_1123,in_1124,in_1125,in_1126,w_44,w_45);
   M50 m23(in_1127,in_1128,in_1129,in_1130,in_1131,in_1132,in_1133,in_1134,in_1135,in_1136,in_1137,in_1138,in_1139,in_1140,in_1141,in_1142,in_1143,in_1144,in_1145,in_1146,in_1147,in_1148,in_1149,in_1150,in_1151,in_1152,in_1153,in_1154,in_1155,in_1156,in_1157,in_1158,in_1159,in_1160,in_1161,in_1162,in_1163,in_1164,in_1165,in_1166,in_1167,in_1168,in_1169,in_1170,in_1171,in_1172,in_1173,in_1174,in_1175,w_46,w_47);
   M50 m24(in_1176,in_1177,in_1178,in_1179,in_1180,in_1181,in_1182,in_1183,in_1184,in_1185,in_1186,in_1187,in_1188,in_1189,in_1190,in_1191,in_1192,in_1193,in_1194,in_1195,in_1196,in_1197,in_1198,in_1199,in_1200,in_1201,in_1202,in_1203,in_1204,in_1205,in_1206,in_1207,in_1208,in_1209,in_1210,in_1211,in_1212,in_1213,in_1214,in_1215,in_1216,in_1217,in_1218,in_1219,in_1220,in_1221,in_1222,in_1223,in_1224,w_48,w_49);
   M50 m25(in_1225,in_1226,in_1227,in_1228,in_1229,in_1230,in_1231,in_1232,in_1233,in_1234,in_1235,in_1236,in_1237,in_1238,in_1239,in_1240,in_1241,in_1242,in_1243,in_1244,in_1245,in_1246,in_1247,in_1248,in_1249,in_1250,in_1251,in_1252,in_1253,in_1254,in_1255,in_1256,in_1257,in_1258,in_1259,in_1260,in_1261,in_1262,in_1263,in_1264,in_1265,in_1266,in_1267,in_1268,in_1269,in_1270,in_1271,in_1272,in_1273,w_50,w_51);
   M50 m26(in_1274,in_1275,in_1276,in_1277,in_1278,in_1279,in_1280,in_1281,in_1282,in_1283,in_1284,in_1285,in_1286,in_1287,in_1288,in_1289,in_1290,in_1291,in_1292,in_1293,in_1294,in_1295,in_1296,in_1297,in_1298,in_1299,in_1300,in_1301,in_1302,in_1303,in_1304,in_1305,in_1306,in_1307,in_1308,in_1309,in_1310,in_1311,in_1312,in_1313,in_1314,in_1315,in_1316,in_1317,in_1318,in_1319,in_1320,in_1321,in_1322,w_52,w_53);
   M50 m27(in_1323,in_1324,in_1325,in_1326,in_1327,in_1328,in_1329,in_1330,in_1331,in_1332,in_1333,in_1334,in_1335,in_1336,in_1337,in_1338,in_1339,in_1340,in_1341,in_1342,in_1343,in_1344,in_1345,in_1346,in_1347,in_1348,in_1349,in_1350,in_1351,in_1352,in_1353,in_1354,in_1355,in_1356,in_1357,in_1358,in_1359,in_1360,in_1361,in_1362,in_1363,in_1364,in_1365,in_1366,in_1367,in_1368,in_1369,in_1370,in_1371,w_54,w_55);
   M50 m28(in_1372,in_1373,in_1374,in_1375,in_1376,in_1377,in_1378,in_1379,in_1380,in_1381,in_1382,in_1383,in_1384,in_1385,in_1386,in_1387,in_1388,in_1389,in_1390,in_1391,in_1392,in_1393,in_1394,in_1395,in_1396,in_1397,in_1398,in_1399,in_1400,in_1401,in_1402,in_1403,in_1404,in_1405,in_1406,in_1407,in_1408,in_1409,in_1410,in_1411,in_1412,in_1413,in_1414,in_1415,in_1416,in_1417,in_1418,in_1419,in_1420,w_56,w_57);
   M50 m29(in_1421,in_1422,in_1423,in_1424,in_1425,in_1426,in_1427,in_1428,in_1429,in_1430,in_1431,in_1432,in_1433,in_1434,in_1435,in_1436,in_1437,in_1438,in_1439,in_1440,in_1441,in_1442,in_1443,in_1444,in_1445,in_1446,in_1447,in_1448,in_1449,in_1450,in_1451,in_1452,in_1453,in_1454,in_1455,in_1456,in_1457,in_1458,in_1459,in_1460,in_1461,in_1462,in_1463,in_1464,in_1465,in_1466,in_1467,in_1468,in_1469,w_58,w_59);
   M50 m30(in_1470,in_1471,in_1472,in_1473,in_1474,in_1475,in_1476,in_1477,in_1478,in_1479,in_1480,in_1481,in_1482,in_1483,in_1484,in_1485,in_1486,in_1487,in_1488,in_1489,in_1490,in_1491,in_1492,in_1493,in_1494,in_1495,in_1496,in_1497,in_1498,in_1499,in_1500,in_1501,in_1502,in_1503,in_1504,in_1505,in_1506,in_1507,in_1508,in_1509,in_1510,in_1511,in_1512,in_1513,in_1514,in_1515,in_1516,in_1517,in_1518,w_60,w_61);
   M50 m31(in_1519,in_1520,in_1521,in_1522,in_1523,in_1524,in_1525,in_1526,in_1527,in_1528,in_1529,in_1530,in_1531,in_1532,in_1533,in_1534,in_1535,in_1536,in_1537,in_1538,in_1539,in_1540,in_1541,in_1542,in_1543,in_1544,in_1545,in_1546,in_1547,in_1548,in_1549,in_1550,in_1551,in_1552,in_1553,in_1554,in_1555,in_1556,in_1557,in_1558,in_1559,in_1560,in_1561,in_1562,in_1563,in_1564,in_1565,in_1566,in_1567,w_62,w_63);
   M50 m32(in_1568,in_1569,in_1570,in_1571,in_1572,in_1573,in_1574,in_1575,in_1576,in_1577,in_1578,in_1579,in_1580,in_1581,in_1582,in_1583,in_1584,in_1585,in_1586,in_1587,in_1588,in_1589,in_1590,in_1591,in_1592,in_1593,in_1594,in_1595,in_1596,in_1597,in_1598,in_1599,in_1600,in_1601,in_1602,in_1603,in_1604,in_1605,in_1606,in_1607,in_1608,in_1609,in_1610,in_1611,in_1612,in_1613,in_1614,in_1615,in_1616,w_64,w_65);
   M50 m33(in_1617,in_1618,in_1619,in_1620,in_1621,in_1622,in_1623,in_1624,in_1625,in_1626,in_1627,in_1628,in_1629,in_1630,in_1631,in_1632,in_1633,in_1634,in_1635,in_1636,in_1637,in_1638,in_1639,in_1640,in_1641,in_1642,in_1643,in_1644,in_1645,in_1646,in_1647,in_1648,in_1649,in_1650,in_1651,in_1652,in_1653,in_1654,in_1655,in_1656,in_1657,in_1658,in_1659,in_1660,in_1661,in_1662,in_1663,in_1664,in_1665,w_66,w_67);
   M50 m34(in_1666,in_1667,in_1668,in_1669,in_1670,in_1671,in_1672,in_1673,in_1674,in_1675,in_1676,in_1677,in_1678,in_1679,in_1680,in_1681,in_1682,in_1683,in_1684,in_1685,in_1686,in_1687,in_1688,in_1689,in_1690,in_1691,in_1692,in_1693,in_1694,in_1695,in_1696,in_1697,in_1698,in_1699,in_1700,in_1701,in_1702,in_1703,in_1704,in_1705,in_1706,in_1707,in_1708,in_1709,in_1710,in_1711,in_1712,in_1713,in_1714,w_68,w_69);
   M50 m35(in_1715,in_1716,in_1717,in_1718,in_1719,in_1720,in_1721,in_1722,in_1723,in_1724,in_1725,in_1726,in_1727,in_1728,in_1729,in_1730,in_1731,in_1732,in_1733,in_1734,in_1735,in_1736,in_1737,in_1738,in_1739,in_1740,in_1741,in_1742,in_1743,in_1744,in_1745,in_1746,in_1747,in_1748,in_1749,in_1750,in_1751,in_1752,in_1753,in_1754,in_1755,in_1756,in_1757,in_1758,in_1759,in_1760,in_1761,in_1762,in_1763,w_70,w_71);
   M50 m36(in_1764,in_1765,in_1766,in_1767,in_1768,in_1769,in_1770,in_1771,in_1772,in_1773,in_1774,in_1775,in_1776,in_1777,in_1778,in_1779,in_1780,in_1781,in_1782,in_1783,in_1784,in_1785,in_1786,in_1787,in_1788,in_1789,in_1790,in_1791,in_1792,in_1793,in_1794,in_1795,in_1796,in_1797,in_1798,in_1799,in_1800,in_1801,in_1802,in_1803,in_1804,in_1805,in_1806,in_1807,in_1808,in_1809,in_1810,in_1811,in_1812,w_72,w_73);
   M50 m37(in_1813,in_1814,in_1815,in_1816,in_1817,in_1818,in_1819,in_1820,in_1821,in_1822,in_1823,in_1824,in_1825,in_1826,in_1827,in_1828,in_1829,in_1830,in_1831,in_1832,in_1833,in_1834,in_1835,in_1836,in_1837,in_1838,in_1839,in_1840,in_1841,in_1842,in_1843,in_1844,in_1845,in_1846,in_1847,in_1848,in_1849,in_1850,in_1851,in_1852,in_1853,in_1854,in_1855,in_1856,in_1857,in_1858,in_1859,in_1860,in_1861,w_74,w_75);
   M50 m38(in_1862,in_1863,in_1864,in_1865,in_1866,in_1867,in_1868,in_1869,in_1870,in_1871,in_1872,in_1873,in_1874,in_1875,in_1876,in_1877,in_1878,in_1879,in_1880,in_1881,in_1882,in_1883,in_1884,in_1885,in_1886,in_1887,in_1888,in_1889,in_1890,in_1891,in_1892,in_1893,in_1894,in_1895,in_1896,in_1897,in_1898,in_1899,in_1900,in_1901,in_1902,in_1903,in_1904,in_1905,in_1906,in_1907,in_1908,in_1909,in_1910,w_76,w_77);
   M50 m39(in_1911,in_1912,in_1913,in_1914,in_1915,in_1916,in_1917,in_1918,in_1919,in_1920,in_1921,in_1922,in_1923,in_1924,in_1925,in_1926,in_1927,in_1928,in_1929,in_1930,in_1931,in_1932,in_1933,in_1934,in_1935,in_1936,in_1937,in_1938,in_1939,in_1940,in_1941,in_1942,in_1943,in_1944,in_1945,in_1946,in_1947,in_1948,in_1949,in_1950,in_1951,in_1952,in_1953,in_1954,in_1955,in_1956,in_1957,in_1958,in_1959,w_78,w_79);
   M50 m40(in_1960,in_1961,in_1962,in_1963,in_1964,in_1965,in_1966,in_1967,in_1968,in_1969,in_1970,in_1971,in_1972,in_1973,in_1974,in_1975,in_1976,in_1977,in_1978,in_1979,in_1980,in_1981,in_1982,in_1983,in_1984,in_1985,in_1986,in_1987,in_1988,in_1989,in_1990,in_1991,in_1992,in_1993,in_1994,in_1995,in_1996,in_1997,in_1998,in_1999,in_2000,in_2001,in_2002,in_2003,in_2004,in_2005,in_2006,in_2007,in_2008,w_80,w_81);
   M50 m41(in_2009,in_2010,in_2011,in_2012,in_2013,in_2014,in_2015,in_2016,in_2017,in_2018,in_2019,in_2020,in_2021,in_2022,in_2023,in_2024,in_2025,in_2026,in_2027,in_2028,in_2029,in_2030,in_2031,in_2032,in_2033,in_2034,in_2035,in_2036,in_2037,in_2038,in_2039,in_2040,in_2041,in_2042,in_2043,in_2044,in_2045,in_2046,in_2047,in_2048,in_2049,in_2050,in_2051,in_2052,in_2053,in_2054,in_2055,in_2056,in_2057,w_82,w_83);
   M50 m42(in_2058,in_2059,in_2060,in_2061,in_2062,in_2063,in_2064,in_2065,in_2066,in_2067,in_2068,in_2069,in_2070,in_2071,in_2072,in_2073,in_2074,in_2075,in_2076,in_2077,in_2078,in_2079,in_2080,in_2081,in_2082,in_2083,in_2084,in_2085,in_2086,in_2087,in_2088,in_2089,in_2090,in_2091,in_2092,in_2093,in_2094,in_2095,in_2096,in_2097,in_2098,in_2099,in_2100,in_2101,in_2102,in_2103,in_2104,in_2105,in_2106,w_84,w_85);
   M50 m43(in_2107,in_2108,in_2109,in_2110,in_2111,in_2112,in_2113,in_2114,in_2115,in_2116,in_2117,in_2118,in_2119,in_2120,in_2121,in_2122,in_2123,in_2124,in_2125,in_2126,in_2127,in_2128,in_2129,in_2130,in_2131,in_2132,in_2133,in_2134,in_2135,in_2136,in_2137,in_2138,in_2139,in_2140,in_2141,in_2142,in_2143,in_2144,in_2145,in_2146,in_2147,in_2148,in_2149,in_2150,in_2151,in_2152,in_2153,in_2154,in_2155,w_86,w_87);
   M50 m44(in_2156,in_2157,in_2158,in_2159,in_2160,in_2161,in_2162,in_2163,in_2164,in_2165,in_2166,in_2167,in_2168,in_2169,in_2170,in_2171,in_2172,in_2173,in_2174,in_2175,in_2176,in_2177,in_2178,in_2179,in_2180,in_2181,in_2182,in_2183,in_2184,in_2185,in_2186,in_2187,in_2188,in_2189,in_2190,in_2191,in_2192,in_2193,in_2194,in_2195,in_2196,in_2197,in_2198,in_2199,in_2200,in_2201,in_2202,in_2203,in_2204,w_88,w_89);
   M50 m45(in_2205,in_2206,in_2207,in_2208,in_2209,in_2210,in_2211,in_2212,in_2213,in_2214,in_2215,in_2216,in_2217,in_2218,in_2219,in_2220,in_2221,in_2222,in_2223,in_2224,in_2225,in_2226,in_2227,in_2228,in_2229,in_2230,in_2231,in_2232,in_2233,in_2234,in_2235,in_2236,in_2237,in_2238,in_2239,in_2240,in_2241,in_2242,in_2243,in_2244,in_2245,in_2246,in_2247,in_2248,in_2249,in_2250,in_2251,in_2252,in_2253,w_90,w_91);
   M50 m46(in_2254,in_2255,in_2256,in_2257,in_2258,in_2259,in_2260,in_2261,in_2262,in_2263,in_2264,in_2265,in_2266,in_2267,in_2268,in_2269,in_2270,in_2271,in_2272,in_2273,in_2274,in_2275,in_2276,in_2277,in_2278,in_2279,in_2280,in_2281,in_2282,in_2283,in_2284,in_2285,in_2286,in_2287,in_2288,in_2289,in_2290,in_2291,in_2292,in_2293,in_2294,in_2295,in_2296,in_2297,in_2298,in_2299,in_2300,in_2301,in_2302,w_92,w_93);
   M50 m47(in_2303,in_2304,in_2305,in_2306,in_2307,in_2308,in_2309,in_2310,in_2311,in_2312,in_2313,in_2314,in_2315,in_2316,in_2317,in_2318,in_2319,in_2320,in_2321,in_2322,in_2323,in_2324,in_2325,in_2326,in_2327,in_2328,in_2329,in_2330,in_2331,in_2332,in_2333,in_2334,in_2335,in_2336,in_2337,in_2338,in_2339,in_2340,in_2341,in_2342,in_2343,in_2344,in_2345,in_2346,in_2347,in_2348,in_2349,in_2350,in_2351,w_94,w_95);
   M50 m48(in_2352,in_2353,in_2354,in_2355,in_2356,in_2357,in_2358,in_2359,in_2360,in_2361,in_2362,in_2363,in_2364,in_2365,in_2366,in_2367,in_2368,in_2369,in_2370,in_2371,in_2372,in_2373,in_2374,in_2375,in_2376,in_2377,in_2378,in_2379,in_2380,in_2381,in_2382,in_2383,in_2384,in_2385,in_2386,in_2387,in_2388,in_2389,in_2390,in_2391,in_2392,in_2393,in_2394,in_2395,in_2396,in_2397,in_2398,in_2399,in_2400,w_96,w_97);
   M50 m49(in_2401,in_2402,in_2403,in_2404,in_2405,in_2406,in_2407,in_2408,in_2409,in_2410,in_2411,in_2412,in_2413,in_2414,in_2415,in_2416,in_2417,in_2418,in_2419,in_2420,in_2421,in_2422,in_2423,in_2424,in_2425,in_2426,in_2427,in_2428,in_2429,in_2430,in_2431,in_2432,in_2433,in_2434,in_2435,in_2436,in_2437,in_2438,in_2439,in_2440,in_2441,in_2442,in_2443,in_2444,in_2445,in_2446,in_2447,in_2448,in_2449,w_98,w_99);

endmodule


module M48 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M49 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M49 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M47 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M48 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M48 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M46 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M47 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M47 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M45 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M46 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M46 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M44 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M45 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M45 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M43 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M44 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M44 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M42 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M43 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M43 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M41 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M42 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M42 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M40 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M41 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M41 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M39 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M40 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M40 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M38 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M39 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M39 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M37 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M38 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M38 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M36 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M37 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M37 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M35 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M36 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M36 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M34 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M35 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M35 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M33 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M34 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M34 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M32 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M33 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M33 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M31 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M32 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M32 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M30 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M31 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M31 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M29 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M30 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M30 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M28 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M29 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M29 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M27 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M28 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M28 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M26 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M27 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M27 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M25 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M26 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M26 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M24 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M25 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M25 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M23 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M24 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M24 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M22 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M23 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M23 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M21 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M22 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M22 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M20 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M21 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M21 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M19 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M20 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M20 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M18 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M19 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M19 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M17 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M18 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M18 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M16 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M17 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M17 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M15 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M16 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M16 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M14 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M15 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M15 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M13 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M14 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M14 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M12 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M13 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M13 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M11 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M12 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M12 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M10 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M11 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M11 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M9 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M10 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M10 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M8 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M9 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M9 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M7 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M8 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M8 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M6 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M7 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M7 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M5 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M6 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M6 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M4 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_5;

   M5 m0(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m1(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m2(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m3(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m4(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m5(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m6(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m7(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m8(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m9(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m10(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m11(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m12(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m13(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m14(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m15(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m16(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m17(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m18(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m19(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m20(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m21(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m22(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m23(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m24(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m25(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m26(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m27(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m28(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m29(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m30(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m31(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m32(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m33(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m34(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m35(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m36(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m37(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m38(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m39(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m40(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m41(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m42(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m43(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m44(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m45(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m46(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m47(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m48(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);
   M5 m49(out_0,out_1,out_2,out_3,out_4,out_5,in_0,in_1,in_2,in_3,in_5,in_5);

endmodule


module M3 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_0;

   M4 m0(in_0,in_1,in_2,in_3,in_4,in_5,w_0,w_1,w_2,w_3,w_4);
   
endmodule


module M2 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_5;

	assign out_0 = w_0 + w_1;
	assign out_1 = w_1 & w_2;
	assign out_2 = w_2 | w_3;
	assign out_3 = w_3 + w_4;
	assign out_4 = w_4 & w_0;

   M3 m0(in_0,in_1,in_2,in_3,in_4,in_5,w_0,w_1,w_2,w_3,w_4);
   
endmodule


module M1 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_6;
	wire [16:0] w_7;
	wire [16:0] w_8;
	wire [16:0] w_9;
	wire [16:0] w_10;
	wire [16:0] w_11;
	wire [16:0] w_12;
	wire [16:0] w_13;
	wire [16:0] w_14;
	wire [16:0] w_15;
	wire [16:0] w_16;
	wire [16:0] w_17;
	wire [16:0] w_18;
	wire [16:0] w_19;

	assign w_15 = w_0 + w_1;
	assign w_16 = w_2 & w_3;
	assign w_17 = w_4 | w_5;
	assign w_18 = w_6 + w_7;
	assign w_19 = w_8 & w_9;
	assign out_0 = w_10 | w_15;
	assign out_1 = w_11 + w_16;
	assign out_2 = w_12 & w_17;
	assign out_3 = w_13 | w_18;
	assign out_4 = w_14 + w_19;
   M2 m0(in_0,in_1,in_2,in_3,in_4,in_5,w_0,w_1,w_2,w_3,w_4);
   M2 m1(in_0,in_1,in_2,in_3,in_4,in_5,w_5,w_6,w_7,w_8,w_9);
   M2 m2(in_0,in_1,in_2,in_3,in_4,in_5,w_10,w_11,w_12,w_13,w_14);
   M2 m3(in_0,in_1,in_2,in_3,in_4,in_5,w_15,w_16,w_17,w_18,w_19);
   
endmodule

module mux2to1(in_0,in_1,in_2,in_3,in_4,in_5,data_out);
input [16:0] in_0;
input [16:0] in_1;
input [16:0] in_2;
input [16:0] in_3;
input [16:0] in_4;
input [16:0] in_5;
output [16:0] data_out;
reg [16:0] data_out;
always @(in_0,in_1,in_2,in_3,in_4,in_5)
	begin
		if(in_5== 0)
			data_out =in_0+in_1+in_2+in_3+in_4+in_5+;
		else
			data_out = in_4 & in_5;

	end
endmodule


module M0 (in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
   input [16:0] in_0;
   input [16:0] in_1;
   input [16:0] in_2;
   input [16:0] in_3;
   input [16:0] in_4;
   input [16:0] in_5;
   output [16:0] out_0;
   output [16:0] out_1;
   output [16:0] out_2;
   output [16:0] out_3;
   output [16:0] out_4;

	wire [16:0] w_0;
	wire [16:0] w_1;
	wire [16:0] w_2;
	wire [16:0] w_3;
	wire [16:0] w_4;
	wire [16:0] w_6;
	wire [16:0] w_7;
	wire [16:0] w_8;
	wire [16:0] w_9;
	wire [16:0] w_10;
	wire [16:0] w_11;
	wire [16:0] w_12;
	wire [16:0] w_13;
	wire [16:0] w_14;
	wire [16:0] w_15;

	assign out_0 =  w_0;
	assign out_1 =  w_1;
	assign out_2 =  w_2;
	assign out_3 =  w_3;
   assign out_4 =  w_4;
	assign w_0 = w_6 & w_11;
	assign w_1 = w_7 | w_12;
	assign w_2 = w_8 + w_13;
	assign w_3 = w_9 & w_14;
	assign w_4 = w_10 | w_15;

   M1 m0(in_0,in_1,in_2,in_3,in_4,in_5,w_6,w_7,w_8,w_9,w_10);
   M1 m1(in_0,in_1,in_2,in_3,in_4,in_5,w_11,w_12,w_13,w_14,w_15);
   mux2to1  m2(in_5,w_0,w_1,w_2,w_3,w_4,out_4);


endmodule
