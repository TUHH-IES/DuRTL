module FiftyModule_tb;
reg [16:0] in_0, in_1, in_2, in_3, in_4, in_5;
output [16:0]out_0,out_1,out_2,out_3,out_4;
M0 test(in_0,in_1,in_2,in_3,in_4,in_5,out_0,out_1,out_2,out_3,out_4);
initial begin
in_0 = 17'b00000000000000000;
in_1 = 17'b00000000000000000;
in_2 = 17'b00000000000000000;
in_3 = 17'b00000000000000000;
in_4 = 17'b00000000000000000;
in_5 = 17'b00000000000000000;
#2
in_0 = 17'b00000000001111111;
in_1 = 17'b00000000011111111;
in_2 = 17'b00000000111111111;
in_3 = 17'b00000001111111111;
in_4 = 17'b00000011111111111;
in_5 = 17'b00000111111111111;
#4
in_0 = 17'b00000000000000000;
in_1 = 17'b00000000000000000;
in_2 = 17'b00000000000000000;
in_3 = 17'b11111111111111111;
in_4 = 17'b00000000000000000;
in_5 = 17'b00000000000000000;
#6
in_0 = 17'b11111111100000000;
in_1 = 17'b11111111000000000;
in_2 = 17'b11111111000000000;
in_3 = 17'b11111111111111111;
in_4 = 17'b11111111000000000;
in_5 = 17'b11111111000000000;
#8
in_0 = 17'b00000000011111111;
in_1 = 17'b00000000011111111;
in_2 = 17'b00000000011111111;
in_3 = 17'b11111111111111111;
in_4 = 17'b00000000011111111;
in_5 = 17'b00000000011111111;
#10
in_0 = 17'b00000000000000000;
in_1 = 17'b00000000000000000;
in_2 = 17'b00000000000000000;
in_3 = 17'b00000000111111110;
in_4 = 17'b00000000000000000;
in_5 = 17'b00000000000000000;
#12
in_0 = 17'b11111111000000000;
in_1 = 17'b11111111100000000;
in_2 = 17'b11111111110000000;
in_3 = 17'b11111111111111111;
in_4 = 17'b11111111111100000;
in_5 = 17'b11111111111110000;
#14
in_0 = 17'b11111111111111110;
in_1 = 17'b11111111111111110;
in_2 = 17'b11111111111111110;
in_3 = 17'b11111111111111110;
in_4 = 17'b11111111111111110;
in_5 = 17'b11111111111111110;
end
initial
begin
	$dumpfile("../../examples/PathMaker/../Fifty/FiftyModule.vcd");
	$dumpvars();
end
endmodule
